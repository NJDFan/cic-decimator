------------------------------------------------------------------------
-- CIC Decimator {{ name }}
--
--  Summary:
--      Stages: {{ stages }}
--      Decimation Ratio: {{ ratio }}
--      Input Data Range: {{ input_min }}-{{ input_max }}
--      Output Data Range: {{ output_min }}-{{ output_max }}
--
--  Usage:
--      Data is accepted on the in_data any time in_valid = '1'.
--      Every {{ ratio }} times the data is input, the out_data is
--      updated and out_valid goes high for one clock.
-- 
--      There is no flow control either in or out; {{ name }} can accept
--      input data on every clock and expects that downstream logic can
--      either process or defer output data on the same clock it is
--      generated.
--
--      Note that out_data will remain stable even after out_valid goes
--      low again; so out_valid can be considered to be a new_data flag
--      rather than a valid.
--
------------------------------------------------------------------------
-- Generated {{ now }}
-- Generated by Rob Gaddi's {{ program }}.
--
-- This file is a generated output product, and is unencumbered by
-- any license restrictions that may appear in the {{ program }}
-- license; see LICENSE.TXT for more details.
------------------------------------------------------------------------

-- This file is expected to appear in library {{ work }} 

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity {{ name }} is
    port (
        in_data     : in  {{ input_dtype }};
        in_valid    : in  std_logic;
        out_data    : out {{ output_dtype }};
        out_valid   : out std_logic;
    
        clk : in std_logic;
        {{ "arst" if async_reset else "rst" }} : in std_logic
    );
end entity {{ name }};

architecture Behavioral of {{ name }} is

    subtype dtype is {{ output_dtype }};
    type dtype_array is array(natural range <>) of dtype;
    subtype ta_dtype  is dtype_array({{stages}} downto 1);
    subtype tex_dtype is dtype_array({{stages}} downto 0);
    
    constant DATA_RESET : ta_dtype := (others => (others => '0'));
    signal integrator : ta_dtype := DATA_RESET;
    signal comb       : ta_dtype := DATA_RESET;
    signal comb_x     : ta_dtype := DATA_RESET;
    
    -- High when a given stage in either the integrator or comb has newly
    -- updated data.
    signal int_flag   : std_logic_vector({{stages}} downto 1) := (others => '0');
    signal comb_flag  : std_logic_vector({{stages}} downto 1) := (others => '0');

    -- High when the next int_flag'high should cause the combs to fire.
    signal decimate_flag : std_logic;

begin

    -- For any CIC filter the integrators run on the fast
    -- side, and the combs run on the slow side.  This being
    -- a decimating filter, that puts the integrators on the
    -- input and the combs on the output.

    INTEGRATORS: process(clk {{", arst" if async_reset}})
        variable d     : dtype;
        variable data  : tex_dtype;
        variable flag  : std_logic_vector({{stages}} downto 0);
    begin
        {% if async_reset %}
        -- Asynchronous reset
        if (arst = '1') then
            int_flag   <= (others => '0');
            integrator <= DATA_RESET;
            
        elsif rising_edge(clk) then
        {% else %}
        if rising_edge(clk) then
        {% endif %}
            -- Update the integrator data
            d := RESIZE(in_data, out_data'length);
            data(integrator'range) := integrator;
            data(0) := d;
            flag := int_flag & in_valid;
            
            for i in integrator'range loop
                if flag(i-1) = '1' then
                    integrator(i) <= data(i) + data(i-1);
                end if;
            end loop;
            
            -- Shift the data valid shift register
            int_flag <= flag(int_flag'high-1 downto 0);
            
            {% if not async_reset %}
            -- Synchronous reset
            if rst = '1' then
                int_flag   <= (others => '0');
                integrator <= DATA_RESET;
            end if;
            {% endif %}
        end if;
    end process INTEGRATORS;
    
    DECIMATION_COUNTER: process(clk {{", arst" if async_reset}})
        variable counter : integer range 0 to {{ratio-1}} := 0;
    begin
        {% if async_reset %}
        -- Asynchronous reset
        if (arst = '1') then
            counter := 0;
            decimate_flag <= '0';
            
        elsif rising_edge(clk) then
        {% else %}
        if rising_edge(clk) then
        {% endif %}
            if int_flag(int_flag'high) = '1' then
                decimate_flag <= '0';
                case counter is
                    when {{ratio - 1}} =>
                        counter := 0;
                    when {{ratio - 2}} =>
                        counter := counter + 1;
                        decimate_flag <= '1';
                    when others =>
                        counter := counter + 1;
                end case;
            end if;
            
            {% if not async_reset %}
            -- Synchronous reset
            if rst = '1' then
                counter := 0;
                decimate_flag <= '0';
            end if;
            {% endif %}
        end if;
    end process DECIMATION_COUNTER;
    
    COMBS: process(clk {{", arst" if async_reset}})
        variable data  : tex_dtype;
        variable flag  : std_logic_vector({{stages}} downto 0);
    begin
        {% if async_reset %}
        -- Asynchronous reset
        if (arst = '1') then
            comb_flag <= (others => '0');
            comb <= DATA_RESET;
            comb_x <= DATA_RESET;
            
        elsif rising_edge(clk) then
        {% else %}
        if rising_edge(clk) then
        {% endif %}
            -- Update the comb data
            data := comb & integrator(integrator'high);
            flag := comb_flag & (int_flag(int_flag'high) and decimate_flag);
            
            for i in comb'range loop
                if flag(i-1) = '1' then
                    comb(i) <= data(i-1) - comb_x(i);
                    comb_x(i) <= data(i-1);
                end if;
            end loop;
            
            -- Shift the data valid shift register
            comb_flag <= flag(comb_flag'high-1 downto 0);
            
            {% if not async_reset %}
            -- Synchronous reset
            if rst = '1' then
                comb_flag <= (others => '0');
                comb <= DATA_RESET;
                comb_x <= DATA_RESET;
            end if;
            {% endif %}
        end if;
    end process COMBS;
    
    out_data  <= comb(comb'high);
    out_valid <= comb_flag(comb_flag'high);

end architecture Behavioral;
