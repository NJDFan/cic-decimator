------------------------------------------------------------------------
-- CIC Decimator {{ name }}
--
--  Summary:
--      Stages: {{ stages }}
--      Decimation Ratio: {{ ratio }}
--      Input Data Range: {{ input_min }}-{{ input_max }}
--      Output Data Range: {{ output_min }}-{{ output_max }}
--
--  Usage:
--      Data is accepted on the in_data any time in_valid = '1'.
--      Every {{ ratio }} times the data is input, the out_data is
--      updated and out_valid goes high for one clock.
-- 
--      There is no flow control either in or out; {{ name }} can accept
--      input data on every clock and expects that downstream logic can
--      either process or defer output data on the same clock it is
--      generated.
--
--      Note that out_data will remain stable even after out_valid goes
--      low again; so out_valid can be considered to be a new_data flag
--      rather than a valid.
--
------------------------------------------------------------------------
-- Generated {{ now }}
-- Generated by Rob Gaddi's {{ program }}.
--
-- This file is a generated output product, and is unencumbered by
-- any license restrictions that may appear in the {{ program }}
-- license; see LICENSE.TXT for more details.
------------------------------------------------------------------------

-- This file is expected to appear in library {{ work }} 

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity {{ name }} is
    port (
        in_data     : in  {{ dtype }}({{ input_bits-1 }} downto 0);
        in_valid    : in  std_logic;
        out_data    : out {{ dtype }}({{ output_bits-1 }} downto 0);
        out_valid   : out std_logic;
    
        clk : in std_logic;
        {{ "arst" if async_reset else "rst" }} : in std_logic
    );
end entity {{ name }};

architecture Behavioral of {{ name }} is

    {% for w in stage_widths %}
    signal data{{ loop.index0 }} : {{ dtype }}({{ w-1 }} downto 0);
    {% endfor %}


    subtype dtype is {{ dtype }}({{ output_bits-1 }} downto 0);
    type dtype_array is array(natural range <>) of dtype;
    subtype ta_dtype  is dtype_array({{stages}} downto 1);
    subtype tex_dtype is dtype_array({{stages}} downto 0);
    
    constant DATA_RESET : ta_dtype := (others => (others => '0'));
    signal integrator : ta_dtype := DATA_RESET;
    signal comb       : ta_dtype := DATA_RESET;
    signal comb_x     : ta_dtype := DATA_RESET;
    
    -- High when a given stage in either the integrator or comb has newly
    -- available data.  Index matches with the stage number; highest is
    -- the output data valid.
    signal stage_flag       : std_logic_vector({{stages*2}} downto 0) := (others => '0');
    signal stage_flag_reg   : std_logic_vector({{stages*2}} downto 1) := (others => '0');
    
    -- High when the next data through the integrators should cause the
    -- combs to fire.
    signal counter : integer range 0 to {{ratio-1}} := 0;
    signal decimate_flag : boolean;

    signal async_r, sync_r : boolean;

    function drop_lsbs(x, ref : {{dtype}}) return {{dtype}} is
    begin
        if x'length < ref'length then
            return RESIZE(x, ref'length);
        else
            return RESIZE(SHIFT_RIGHT(x, x'length-ref'length), ref'length);
        end if;
    end function drop_lsbs;

begin

    -- Reset conditioning
    {% if async_reset %}
    async_r <= (arst = '1');
    sync_r  <= false;
    {% else %}
    async_r <= false;
    sync_r  <= (rst = '1');
    {% endif %}

    -- Walk a data ready flag through the stages
    SHIFT_FLAG: process(clk, async_r)
    begin
        if async_r then
            stage_flag_reg <= (others => '0');
        elsif rising_edge(clk) then
            stage_flag_reg <= stage_flag({{stages*2-1}} downto 0);
            
            -- Comb flags only set when the decimator allows it
            if not decimate_flag then
                stage_flag_reg({{stages}}) <= '0';
            end if;
            
            if sync_r then
                stage_flag_reg <= (others => '0');
            end if;
        end if;
    end process SHIFT_FLAG;

    -- For any CIC filter the integrators run on the fast
    -- side, and the combs run on the slow side.  This being
    -- a decimating filter, that puts the integrators on the
    -- input and the combs on the output.
    
    -----------------------------------------------------------------------
    --  Integrators
    -----------------------------------------------------------------------
    
    {% for i in range(stages) %}
    
    INTEGRATOR{{ i }}: process(clk, async_r)
    begin
        if async_r then
            data{{i}} <= (others => '0');
        elsif rising_edge(clk) then
            if (stage_flag({{i}}) = '1') then
            {% if i == 0 %}
                data{{i}} <= data{{i}} + drop_lsbs(in_data, data{{i}});
            {% else %}
                data{{i}} <= data{{i}} + drop_lsbs(data{{i-1}}, data{{i}});
            {% endif %}
            end if;
            if sync_r then
                data{{i}} <= (others => '0');
            end if;
        end if;
    end process INTEGRATOR{{ i }};
        
    {% endfor %}

    -----------------------------------------------------------------------
    --  Decimation
    -----------------------------------------------------------------------
    
    DECIMATION_COUNTER: process(clk, async_r)
        variable counter : integer range 0 to {{ratio-1}} := 0;
    begin
        if async_r then
            counter <= 0;
            
        elsif rising_edge(clk) then
            if stage_flag({stages-1}) = '1' then
                if decimate_flag then
                    counter <= 0;
                else
                    counter <= counter + 1;
                end if;
            end if;
            
            if sync_r then
                counter <= 0;
            end if;
        end if;
    end process DECIMATION_COUNTER;
    
    decimate_flag <= (counter = {{ratio-1}});
    
    -----------------------------------------------------------------------
    --  Combs
    -----------------------------------------------------------------------
    
    {% for i in range(stages, stages*2) %}
    
    COMB{{i}}: process(clk, async_r)
        variable last : {{dtype}}(data{{i}}'range); 
    begin
        if async_r then
            last := (others => '0');
            data{{i}} <= (others => '0');
            
        elsif rising_edge(clk) then
            if (stage_flag({{i}}) = '1') then
                data{{i}} <= drop_lsbs(data{{i-1}}, last) - last;
                last := drop_lsbs(data{{i-1}}, last);
            end if;
            
            if sync_r then
                last := (others => '0');
                data{{i}} <= (others => '0');
            end if;
        end if;
    end process COMB{{i}};
        
    {% endfor %}
    
    -- Final data truncation
    data{{stages*2}} <= drop_lsbs(data{{stages*2-1}}, data{{stages*2}});
    
    -----------------------------------------------------------------------
    --  Data outputs
    -----------------------------------------------------------------------
    
    out_data  <= data{{stages*2}};
    out_valid <= stage_flag({{stages*2}});

end architecture Behavioral;
